

module mfp_register_r
#(
    parameter WIDTH = 32
)
(
    input                        clk,
    input                        rst,
    input      [ WIDTH - 1 : 0 ] d,
    input                        wr,
    output reg [ WIDTH - 1 : 0 ] q
);
    always @ (posedge clk)
        if(~rst)
            q <= { WIDTH { 1'b0 } };
        else
            if(wr) q <= d;
endmodule